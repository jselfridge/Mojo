
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//
// control.v
// Implements the control law within the avionics board.
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//

module control
  (

  // Clock and reset
  input clk,
  input rst,

  // Command input signals
  //input [7:0] radio_sig,
  //input ch1_isig,
  //input ch2_isig,
  //input ch3_isig,
  //input ch4_isig,
  //input ch5_isig,
  //input ch6_isig,
  //input ch7_isig,

  // Command input values
  //output [9:0] radio_val [7:0],
  //output [9:0] ch1_ival,
  //output [9:0] ch2_ival,
  //output [9:0] ch3_ival,
  //output [9:0] ch4_ival,
  //output [9:0] ch5_ival,
  //output [9:0] ch6_ival,
  //output [9:0] ch7_ival

  );




endmodule



