
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//
// spi_slave_tb.v
// Test bench for the 'spi_slave' module.
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//

module spi_slave_tb ();

  // Assign test stimulus at certain points
  initial begin

    $finish;

  end

endmodule



