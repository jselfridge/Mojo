
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//
// bcd2ascii_tb.v
// Test bench for the 'bcd2ascii' module.
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//

module bcd2ascii_tb ();

  // Number of digits in BCD representation
  localparam BDC_LEN = 3;

  // Test bench inputs
  reg [(4*BCD_LEN)-1:0] bcd;

  // Test bench outputs
  //wire [(8*BCD_LEN)-1:0] ascii;

  // Assign test stimulus at certain points
  initial begin

    bcd = 12'b0000_0000_0000;  #10;  // 000
    bcd = 12'b0000_0000_0001;  #10;  // 001
    bcd = 12'b0000_0000_0100;  #10;  // 004
    bcd = 12'b0000_0000_0111;  #10;  // 007
    bcd = 12'b0000_0000_1001;  #10;  // 009

    bcd = 12'b0000_0010_0000;  #10;  // 020
    bcd = 12'b0000_0010_0001;  #10;  // 021
    bcd = 12'b0000_0010_0100;  #10;  // 024
    bcd = 12'b0000_0010_0111;  #10;  // 027
    bcd = 12'b0000_0010_1001;  #10;  // 029

    bcd = 12'b0000_1001_0000;  #10;  // 090
    bcd = 12'b0000_1001_0001;  #10;  // 091
    bcd = 12'b0000_1001_0100;  #10;  // 094
    bcd = 12'b0000_1001_0111;  #10;  // 097
    bcd = 12'b0000_1001_1001;  #10;  // 099

    bcd = 12'b0011_0000_0000;  #10;  // 300
    bcd = 12'b0011_0000_0001;  #10;  // 301
    bcd = 12'b0011_0000_0100;  #10;  // 304
    bcd = 12'b0011_0000_0111;  #10;  // 307
    bcd = 12'b0011_0000_1001;  #10;  // 309

    bcd = 12'b1001_0000_0000;  #10;  // 900
    bcd = 12'b1001_0000_0001;  #10;  // 901
    bcd = 12'b1001_0000_0100;  #10;  // 904
    bcd = 12'b1001_0000_0111;  #10;  // 907
    bcd = 12'b1001_0000_1001;  #10;  // 909

    bcd = 12'b0110_0101_0000;  #10;  // 650
    bcd = 12'b0110_0101_0001;  #10;  // 651
    bcd = 12'b0110_0101_0100;  #10;  // 654
    bcd = 12'b0110_0101_0111;  #10;  // 657
    bcd = 12'b0110_0101_1001;  #10;  // 659

    $finish;

  end

endmodule



