
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//
// bcd2ascii_tb.v
// Test bench for the 'bcd2ascii' module.
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~//

module bcd2ascii_tb ();

  // Number of characters in number representation
  localparam CHAR_LEN = 2'd3;

  // Test bench inputs
  reg [(4*CHAR_LEN)-1:0] bcd;

  // Test bench outputs
  wire [(8*CHAR_LEN)-1:0] ascii;

  // Connect 'bcd2ascii' module
  bcd2ascii #(
    .CHAR_LEN(3) )
    DUT_bcd2ascii (
    .bcd(bcd),
    .ascii(ascii) );

  // Assign test stimulus at certain points
  initial begin

    bcd = 12'b0000_0000_0000;  #100;  // 000
    bcd = 12'b0000_0000_0001;  #100;  // 001
    bcd = 12'b0000_0000_0100;  #100;  // 004
    bcd = 12'b0000_0000_0111;  #100;  // 007
    bcd = 12'b0000_0000_1001;  #100;  // 009

    bcd = 12'b0000_0010_0000;  #100;  // 020
    bcd = 12'b0000_0010_0001;  #100;  // 021
    bcd = 12'b0000_0010_0100;  #100;  // 024
    bcd = 12'b0000_0010_0111;  #100;  // 027
    bcd = 12'b0000_0010_1001;  #100;  // 029

    bcd = 12'b0000_1001_0000;  #100;  // 090
    bcd = 12'b0000_1001_0001;  #100;  // 091
    bcd = 12'b0000_1001_0100;  #100;  // 094
    bcd = 12'b0000_1001_0111;  #100;  // 097
    bcd = 12'b0000_1001_1001;  #100;  // 099

    bcd = 12'b0011_0000_0000;  #100;  // 300
    bcd = 12'b0011_0000_0001;  #100;  // 301
    bcd = 12'b0011_0000_0100;  #100;  // 304
    bcd = 12'b0011_0000_0111;  #100;  // 307
    bcd = 12'b0011_0000_1001;  #100;  // 309

    bcd = 12'b1001_0000_0000;  #100;  // 900
    bcd = 12'b1001_0000_0001;  #100;  // 901
    bcd = 12'b1001_0000_0100;  #100;  // 904
    bcd = 12'b1001_0000_0111;  #100;  // 907
    bcd = 12'b1001_0000_1001;  #100;  // 909

    bcd = 12'b0110_0101_0000;  #100;  // 650
    bcd = 12'b0110_0101_0001;  #100;  // 651
    bcd = 12'b0110_0101_0100;  #100;  // 654
    bcd = 12'b0110_0101_0111;  #100;  // 657
    bcd = 12'b0110_0101_1001;  #100;  // 659

    bcd = 12'b0000_0000_0000;  #100;  // 000
    #300 $finish;

  end

endmodule



